
package gf_mult_pkg;

    typedef enum logic      {IDLE         = 0,
                             PENDING      = 1} status_e;
endpackage : gf_mult_pkg
