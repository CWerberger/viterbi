
package viterbi_top_pkg;

    typedef enum logic      {IDLE         = 0,
                             PENDING      = 1} status_e;
endpackage : viterbi_top_pkg
